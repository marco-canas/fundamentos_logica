��  CCircuit��  CSerializeHack           ��  CPart              ���  CBuzzer�� 	 CTerminal  ����                           
�  �<�Q                             |��<         ��  6 `  �� 	 CFilament��  CDummyValue  xpxp    1W            �?      �? W 
�  hp}q                           
�  �p�q                            |��           ��`   �� 
 CBattery9V�  � `� `    9V            "@      �? V 
�  � P� e                           
�  � P� e              "@            � d� �         ��   �  ��  CSPDT��  CToggle  *���        
�  8�9�             "@          
�  X�Y�                          
�  x�y�               �            *���         ����P    ��  "� �       
�  0D1Y             "@          
�  PDQY             "@          
�  pDqY               �            "�D     !   ����P                  ���  CWire  (�)�       %�  (p)�       %�  (�q�      %�  p q�       %�   q      %�   	!       %�  X 	!      %�  X�Y!       %�  PXQ�       %��� 
 CCrossOver  �|��        ��Q�      %�  ���       %�0�  �|��        �X�       %�  � �      %�  �X1Y      %�  � � Q       %�  8�9       %�  � 9      %�  x���      %�  �P��       %�  �P�Q      %�  �P�Y       %�  pX�Y      %�  �P�Q       %�  `P�Q       %�  �P�a        %�  H`�a       %�  HPIa        %�  � PIQ       %�  `8aQ        %�  `8i9       %�  hpi9        %�  ��)�      %�  �p)q                    �                             H    ?  G    I  D   7    8   -   : ! ! 6 " " . # # > ' H I ( & ) * ( + ) * , - +  , " / / 4 2 . 5 / 3 1 6 9 7 2 3 ! 5   9 3 8  ; < : = ; < > # = @  E A ? B C A D B  C F @ E G  F  &  '            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 