��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CInverter�� 	 CTerminal  H�]�              @          
�  t���               �            \�t�           ��    ��  CAND
�  ����              @          
�  ����               �          
�  ���               �            �|��           ��    ��  CLogicIn�� 	 CLatchKey  � �� �        
�  ��              @            � ��        ����     ��  � i� w        
�  pq              @            � lt        ����                   ���  CWire  ����       �  ����      �  �I�      �  �p��       �  p�q                    �                                                                          �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 