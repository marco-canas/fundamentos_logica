��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CInverter�� 	 CTerminal  �(�)                          
�  �(�)              @            ��4           ��    �
�  ����     
         @          
�  ����               �            ����           ��    ��  CLogicIn�� 	 CLatchKey  p 	�         
�  � �      
         @            � �         ����     ��  p � '         
�  �  � !                            � � $         ����     ���  CExplode              333333�?�������? A
�   ��      	        �         
�  ,�A�      	        �           �,�           ��    ��  CSchmitt�              333333�?�������? A
�   ��      	        �         
�  ,�A�      	        �           �,�            ��    �� 	 CLogicOut
�  0�E�              @            DxT�     $     ��    ��  COR
�  �x�y     	          �          
�  ����              @          
�  ����              @            �t��     '      ��    ��  CAND
�  ����              @          
�  ����     
         @          
�  ��	�              @            ����     ,      ��    *�
�  �P�Q                          
�  �`�a               �          
�  �X	Y     	          �            �L�d     0      ��                  ���  CWire  XY�      
 4�  X�Y      
 4�  X���     
 4�  � � � !       4�  �  � )       4�  � (�)      4�  �  � !      4�  ����     
 4�  ����      
 4�  ����     
 4�  ����      
 4�  X���     
 4�  � Y     
 4�  p���      4��� 
 CCrossOver  n\td        p(q�       4�  �(q)      4�D�  n\td        �`�a      4�  ��1�      4�  ����       4�  ���      4�  �X�y      	 4�  X�Y     	 4�  �`��       4�  �� �Q       4�  � � ��       4�  @�A�                     �                             :    F  7    N   A   ;       Q       ! ! Q $ I $ ' L ' ( J ( ) ) I , B , - < - . . K 0 O 0 1 G 1 2 2 M A @ 7 5 6  P ; 8 : 9   9 = - < > ? = > @ 5 ?  6 C , C H F B  C G E N 1 ) $ ( K . J M ' 2 L G  P 0 8 O  !             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 